//LABORATORIO 8
//ELECTRONICA DIGITAL I
//GABRIEL ALEXANDER FONG PENAGOS 19722
//TESTBENCH

module testbench();
  reg clk, reset1, enable,loads; //VARIABLES DE ENTRADA DE UN BIT DEL MODULO CONTADOR
  reg [11:0]LOAD; //VALOR DEL LOAD DE 12 BITS QUE LE COLOCAMOS COMO FIJO A LA SALIDA DEL CONTADOR
  wire [11:0]CB; //SALIDA DEL CONTADOR DE 12 BITS

  reg [11:0]Addres; //VARIABLE DE ENTRADA DE 12 BITS PARA EL MODULO ROM
  wire [7:0]DATO;// VARIABLE DE SALIDA DE 7 BITS PARA EL MODULO ROM

  reg [3:0]A,B; //VARIABLE DE ENTRADA PARA EL MODULO ALUU
  reg [2:0]SEL; //VARIABLE DE SELECCION DE LA ALUU
  wire [3:0]OUT;//SALIDA DE LA ALU DE 4 BITS


  contador U1(clk, reset1, enable,loads, LOAD, CB);//MODULO EJERCICIO 1
  ROM U2(Addres, DATO);//MODULO EJERCICIO 2
  ALUU U3(A, B, SEL, OUT);//MODULO EJERCIO 3

  always begin //REALIZAMOS EL RELOJ Y QUE CAMBIE CADA UNIDAD DE TIEMPO
    clk <= 1; #1 clk <= ~clk; #1;
  end


  //REALIZAMOS LAS PRUEBAS DEL MODULO CONTADOR
  initial begin
  reset1 = 1;loads = 0; LOAD = 12'b000000000000; //RESETEAMOS Y LA SEÑAL DEL LOAD APAGADA LE ASIGNAMOS
  #1
  $display("\n");
  $display(" CONTADOR 12 BITS ");
  $display("C \t  R \t E  \t L\t LOAD\t      |\tOUT");
  $monitor("%b \t %b\t %b \t %b \t %b | %b ", clk, reset1, enable,loads, LOAD, CB );
  #1 enable = 1; reset1 = 0; //HABILITAMOS EL ENABLE PARA QUE COMIENCE A CONTAR
  #5 enable = 0;//DESHABILITAMOS ENABLE Y DEJA DE CONTAR
  #3 loads = 1; LOAD = 12'b101010101010; //ENCENDEMOS LA BANDERA DE LOAD Y LE SELECCIONAMOS UN VALOR
  #2 enable = 1;//HABILITAMOS EL ENABLE PARA QUE CUENTE, PERO COMO LOAD SIGUE ENCENDIDO NO CAMBIARA EL VALOR DE SALIDA
  #4 loads = 0;//APAGAMOS LA BANDERA DE LOAD Y SIGUE CONTANDO EN EL VALOR COLOCADO DE LOAD
  #4 loads = 1; LOAD = 12'b101010100000;//VOLVEMOS A HABILITAR LA SEÑAL DE LOAD PERO CON EL ENABLE ENCENDIDO, LOAD TIENE PRIORIDAD SOBRE ENABLE
  #4 loads = 0;//DESHABILITAMOS LA BANDERA DE LOAD Y SIGUE CONTANDO
  #2 enable = 0;// DESHABILITAMOS ENABLE DEJA DE CONTAR
  #1 reset1 = 1;
  end
  //REALIZAMOS LAS PRUEBAS DEL MODULO ROM EN DONDE COLOCAMOS LOS VALORES DEL ADDRESS Y NOS MUESTRA SU VALOR
  initial begin
  #30
  $display("\n");
  $display(" ROM ");
  $display("CLK \t  Addres \t  Dato ");
  $monitor("%b \t %b\t %b ", clk, Addres, DATO);
  Addres = 12'b000000000000;// DIRECCION1 8h00
  #1 Addres = 12'b000000000001; //DIRECCION 2 8h01
  #1 Addres = 12'b000000000010; //DIRECCION 3 8h02
  #1 Addres = 12'b000000000011; //DIRECCION 4 8h03
  #1 Addres = 12'b000000000100; //DIRECCION 5 8h04
  #1 Addres = 12'b000000000111; //DIRECCION 6 8h07
  #1 Addres = 12'b000000001010; //DIRECCION 7 8h10
  #1 Addres = 12'b000000000001; //DIRECCION 8 8h01
  #1 Addres = 12'b000000001000; //DIRECCION 9 8h08
  #1 Addres = 12'b000000010000; //DIRECCION 10 8h16
  #1 Addres = 12'b000000001101; //DIRECCION 11 8h13

  end


//REALIZAMOS LAS PRUEBAS DEL MODULO ALUU Y PROBAMOS TODAS LAS FUNCIONES
  initial begin
  #41
  $display("\n");
  $display(" ALU ");
  $display("CLK \t  A \t B  \t  SEL \tOUT");
  $monitor("%b \t %b\t %b \t %b | %b ", clk, A, B, SEL, OUT );
  A = 4'b1010; B = 4'b0011; SEL = 3'b000; //FUNCION  A AND B
  #1 SEL = 3'b001; //FUNCION A OR B
  #1 SEL = 3'b010; //FUNCION A ADD B
  #1 SEL = 3'b010;//FUNCION A ADD B
  #1 SEL = 3'b011;//ESTA FUNCION NO HACE NADA, COLOCAMOS TODOO el MISMO VALOR DE ANTES
  #1 SEL = 3'b100;//FUNCION A AND ~B
  #1 SEL = 3'b101;//FUNCION A OR ~B
  #1 SEL = 3'b110;//FUNCION A LESS B
  #1 SEL = 3'b111;//FUNCION STL
  #1 A = 4'b010; B = 4'b0011;//POR DEFAULT QUE COLOQUE TODP EN 0
  #2 $finish;
  end

  initial begin                                                                 //INICIAMOS PARA COLOCAR LOS DATOS EN GTK WAVE
        $dumpfile("LAB8_tb.vcd");
        $dumpvars(0, testbench);
      end

endmodule
